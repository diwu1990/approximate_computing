// `include "param_def_8bit_075.sv"
// `include "param_def_8bit_05.sv"
// `include "param_def_8bit_025.sv"
// `include "param_def_8bit_uniform.sv"
// `include "param_def_12bit_uniform.sv"
`include "param_def_16bit_uniform.sv"

